module not_5b (a, o);
  input [4:0] a;
  output [4:0] o;
  
  assign o = ~a;
  
endmodule
